module ha(a,b,sum,c);
input a,b;
output sum,c;
xor g1(sum,a,b);
and g2(c,a,b);
endmodule
module bitmultiplier(a,b,c);
input [1:0]a,b;
output[3:0]c;
wire w1;
and g1(c[0],b[0],a[0]);
ha ha1(a[0]&b[1],a[1]&b[0],c[1],w1);
ha ha2(a[1] &b[1],w1,c[2],c[3]);
endmodule
